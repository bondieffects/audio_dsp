-- LIBRARIES and PACKAGES for i2s_clocks_TB
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity i2s_clocks_TB is
end entity;

-- 5.7 Overview of Simulation Test Benches p. 162
-- 8.4 Test Benches p. 272
architecture i2s_clocks_TB_arch of i2s_clocks_TB is

    -- From I2S Specification:
    -- The system master clock (MCLK) is typically 256 × fS.
    -- The bit clock (SCK) is typically 64 × fS in systems with two
    -- 32-bit words per audio sample. Other word lengths scale SCK accordingly.
    constant MCLK_HALF_PERIOD : time := 40.69 ns; -- half period for 12.288MHz clock (1/(12.288MHz*2))
    constant WS_PERIOD : time := 20833.33 ns;     -- 12.288MHz / 256 = 48kHz  
    constant BCLK_PERIOD : time := 651.04 ns;     -- 12.288MHz / 8 = 1.536MHz

    -- Component declaration for DUT
    component i2s_clocks
        port (
            -- Inputs
            i2s_mclk : in std_logic;        -- 12.288MHz master clock from audio_pll
            reset_n : in std_logic;         -- Active low reset

            -- Outputs
            i2s_bclk : out std_logic;       -- 1.536MHz bit clock
            i2s_ws : out std_logic          -- 48kHz word select clock
        );
    end component;

    -- Signal declarations
    signal i2s_mclk_TB : std_logic := '0';  -- 12.288MHz master clock
    signal reset_n_TB : std_logic := '0';   -- Active low reset
    signal i2s_bclk_TB : std_logic;         -- 1.536MHz bit clock
    signal i2s_ws_TB : std_logic;           -- 48kHz word select clock

begin

    -- DUT instantiation
    DUT1: i2s_clocks
        port map (
            i2s_mclk => i2s_mclk_TB,
            reset_n => reset_n_TB,
            i2s_bclk => i2s_bclk_TB,
            i2s_ws => i2s_ws_TB
        );


    -- Free-running 12.288 MHz master clock from
    -- https://www.embeddedrelated.com/showarticle/266/vhdl-tutorial-combining-clocked-and-sequential-logic.php
    i2s_mclk_proc : process
    begin
        i2s_mclk_TB <= '0';
        wait for MCLK_HALF_PERIOD;
        i2s_mclk_TB <= '1';
        wait for MCLK_HALF_PERIOD;
    end process;

    -- Reset stimulus process
    stim_proc : process
    begin
        reset_n_TB <= '0';
        wait for 200 ns;
        reset_n_TB <= '1';
        wait;                     -- hold forever
    end process;

    -- Simple monitoring process (no automated checks to avoid ModelSim issues)
    MONITOR: process
    begin
        -- Wait for reset release
        wait until reset_n_TB = '1';
        report "Reset released - monitoring started" severity note;

        -- Just wait and let the simulation run
        wait for 3 * WS_PERIOD;  -- Run long enough to see multiple WS cycles
        report "Monitoring complete - check waveforms manually" severity note;
        report "Expected BCLK period: 651.04ns (1.536MHz)" severity note;
        report "Expected WS period: 20833.33ns (48kHz)" severity note;
        
        report "TB finished" severity failure;  -- Stop simulation cleanly
    end process;

end architecture i2s_clocks_TB_arch;